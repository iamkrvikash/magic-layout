* SPICE3 file created from inverter.ext - technology: scmos

.option scale=0.2u

M1000 a_7_n19# a_1_n12# IN IN nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 a_7_n19# a_1_n12# VDD VDD pfet w=8 l=2
+  ad=40 pd=26 as=40 ps=26
C0 VDD IN 2.38fF
