magic
tech scmos
timestamp 1604044583
<< nwell >>
rect 0 -12 45 12
<< pwell >>
rect 0 -51 45 -12
<< ntransistor >>
rect 12 -29 14 -21
rect 31 -29 33 -21
rect 15 -36 19 -34
rect 26 -36 30 -34
<< ptransistor >>
rect 11 -4 15 -1
rect 30 -4 34 -1
<< ndiffusion >>
rect 7 -25 12 -21
rect 10 -29 12 -25
rect 14 -22 19 -21
rect 14 -26 15 -22
rect 14 -29 19 -26
rect 15 -34 19 -29
rect 26 -22 31 -21
rect 30 -26 31 -22
rect 26 -29 31 -26
rect 33 -25 38 -21
rect 33 -29 35 -25
rect 26 -34 30 -29
rect 15 -37 19 -36
rect 26 -37 30 -36
<< pdiffusion >>
rect 10 -4 11 -1
rect 15 -4 16 -1
rect 29 -4 30 -1
rect 34 -4 35 -1
<< ndcontact >>
rect 6 -29 10 -25
rect 15 -26 19 -22
rect 26 -26 30 -22
rect 35 -29 39 -25
rect 15 -41 19 -37
rect 26 -41 30 -37
<< pdcontact >>
rect 6 -4 10 0
rect 16 -4 20 0
rect 25 -4 29 0
rect 35 -4 39 0
<< psubstratepcontact >>
rect 6 -48 10 -44
rect 35 -48 39 -44
<< nsubstratencontact >>
rect 6 5 10 9
rect 35 5 39 9
<< polysilicon >>
rect 11 -1 15 1
rect 30 -1 34 1
rect 11 -6 15 -4
rect 30 -6 34 -4
rect 12 -17 14 -6
rect 31 -10 33 -6
rect 21 -12 33 -10
rect 12 -19 24 -17
rect 12 -21 14 -19
rect 31 -21 33 -12
rect 12 -31 14 -29
rect 31 -31 33 -29
rect 13 -36 15 -34
rect 19 -36 26 -34
rect 30 -36 34 -34
<< polycontact >>
rect 17 -13 21 -9
rect 24 -19 28 -15
rect 21 -34 25 -30
<< metal1 >>
rect 10 5 35 9
rect 6 0 9 5
rect 36 0 39 5
rect 16 -9 19 -4
rect 16 -13 17 -9
rect 16 -22 19 -13
rect 26 -15 29 -4
rect 28 -19 29 -15
rect 26 -22 29 -19
rect 6 -44 9 -29
rect 36 -44 39 -29
rect 10 -48 35 -44
<< labels >>
rlabel metal1 19 7 19 7 5 VDD
rlabel metal1 19 -46 19 -46 1 GND
rlabel polycontact 19 -10 19 -10 1 Q
rlabel polycontact 26 -17 26 -17 1 Q_Bar
rlabel polycontact 22 -32 22 -32 1 WL
rlabel ndcontact 16 -40 16 -40 1 BL
rlabel ndcontact 27 -40 27 -40 1 BLB
<< end >>
